LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY FULLADDER_g2 IS PORT(A        : in  STD_LOGIC;
      			 B        : in  STD_LOGIC;
      			 CARRY_IN : in  STD_LOGIC;
      			 SUM      : out STD_LOGIC;
      			 CARRY    : out STD_LOGIC);
END FULLADDER_g2;

ARCHITECTURE STRUCTURAL of FULLADDER_g2 is
COMPONENT ORGATE  PORT (X : in  STD_LOGIC;
		       Y : in  STD_LOGIC;
		       Z : out STD_LOGIC);
END COMPONENT;

COMPONENT HALFADDER PORT (U    : in  STD_LOGIC;
      			  V    : in  STD_LOGIC;
      			  SUM  : out STD_LOGIC;
      			  CARRY: out STD_LOGIC);
END COMPONENT;

 SIGNAL�W_SUM   : STD_LOGIC;�
 SIGNAL�W_CARRY1: STD_LOGIC;
 SIGNAL�W_CARRY2: STD_LOGIC;
BEGIN
MODULE1: HALFADDER PORT MAP (A,B,W_SUM,W_CARRY1);
MODULE2: HALFADDER PORT MAP (W_SUM,CARRY_IN,SUM,W_CARRY2);
MODULE3: ORGATE    PORT MAP (W_CARRY1,W_CARRY2,CARRY);
END STRUCTURAL;

