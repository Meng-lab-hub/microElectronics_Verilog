LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY HALFADDER IS 
 PORT(U,V:         IN  STD_LOGIC; 
      SUM, CARRY : OUT STD_LOGIC); 
END HALFADDER; 

ARCHITECTURE RTL_HALFADDER OF HALFADDER IS 
BEGIN 
  SUM 	<= U XOR V; 
  CARRY <= U AND V;
END; 
